// system.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_clk,                 //             clk.clk
		output wire        hps_0_h2f_reset_reset_n, // hps_0_h2f_reset.reset_n
		output wire [14:0] memory_mem_a,            //          memory.mem_a
		output wire [2:0]  memory_mem_ba,           //                .mem_ba
		output wire        memory_mem_ck,           //                .mem_ck
		output wire        memory_mem_ck_n,         //                .mem_ck_n
		output wire        memory_mem_cke,          //                .mem_cke
		output wire        memory_mem_cs_n,         //                .mem_cs_n
		output wire        memory_mem_ras_n,        //                .mem_ras_n
		output wire        memory_mem_cas_n,        //                .mem_cas_n
		output wire        memory_mem_we_n,         //                .mem_we_n
		output wire        memory_mem_reset_n,      //                .mem_reset_n
		inout  wire [31:0] memory_mem_dq,           //                .mem_dq
		inout  wire [3:0]  memory_mem_dqs,          //                .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,        //                .mem_dqs_n
		output wire        memory_mem_odt,          //                .mem_odt
		output wire [3:0]  memory_mem_dm,           //                .mem_dm
		input  wire        memory_oct_rzqin,        //                .oct_rzqin
		output wire [7:0]  pwm_input_0_export,      //     pwm_input_0.export
		input  wire        reset_reset_n            //           reset.reset_n
	);

	wire         mm_bridge_0_m0_waitrequest;            // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [7:0] mm_bridge_0_m0_readdata;               // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;            // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire   [3:0] mm_bridge_0_m0_address;                // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                   // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire   [0:0] mm_bridge_0_m0_byteenable;             // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;          // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire   [7:0] mm_bridge_0_m0_writedata;              // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                  // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;             // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire         mm_interconnect_0_pio_0_s1_chipselect; // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;   // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;    // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;      // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;  // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         rst_controller_reset_out_reset;        // rst_controller:reset_out -> [mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, pio_0:reset_n]

	system_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (2)
	) hps_0 (
		.mem_a       (memory_mem_a),            //         memory.mem_a
		.mem_ba      (memory_mem_ba),           //               .mem_ba
		.mem_ck      (memory_mem_ck),           //               .mem_ck
		.mem_ck_n    (memory_mem_ck_n),         //               .mem_ck_n
		.mem_cke     (memory_mem_cke),          //               .mem_cke
		.mem_cs_n    (memory_mem_cs_n),         //               .mem_cs_n
		.mem_ras_n   (memory_mem_ras_n),        //               .mem_ras_n
		.mem_cas_n   (memory_mem_cas_n),        //               .mem_cas_n
		.mem_we_n    (memory_mem_we_n),         //               .mem_we_n
		.mem_reset_n (memory_mem_reset_n),      //               .mem_reset_n
		.mem_dq      (memory_mem_dq),           //               .mem_dq
		.mem_dqs     (memory_mem_dqs),          //               .mem_dqs
		.mem_dqs_n   (memory_mem_dqs_n),        //               .mem_dqs_n
		.mem_odt     (memory_mem_odt),          //               .mem_odt
		.mem_dm      (memory_mem_dm),           //               .mem_dm
		.oct_rzqin   (memory_oct_rzqin),        //               .oct_rzqin
		.h2f_rst_n   (hps_0_h2f_reset_reset_n), //      h2f_reset.reset_n
		.h2f_axi_clk (clk_clk),                 //  h2f_axi_clock.clk
		.h2f_AWID    (),                        // h2f_axi_master.awid
		.h2f_AWADDR  (),                        //               .awaddr
		.h2f_AWLEN   (),                        //               .awlen
		.h2f_AWSIZE  (),                        //               .awsize
		.h2f_AWBURST (),                        //               .awburst
		.h2f_AWLOCK  (),                        //               .awlock
		.h2f_AWCACHE (),                        //               .awcache
		.h2f_AWPROT  (),                        //               .awprot
		.h2f_AWVALID (),                        //               .awvalid
		.h2f_AWREADY (),                        //               .awready
		.h2f_WID     (),                        //               .wid
		.h2f_WDATA   (),                        //               .wdata
		.h2f_WSTRB   (),                        //               .wstrb
		.h2f_WLAST   (),                        //               .wlast
		.h2f_WVALID  (),                        //               .wvalid
		.h2f_WREADY  (),                        //               .wready
		.h2f_BID     (),                        //               .bid
		.h2f_BRESP   (),                        //               .bresp
		.h2f_BVALID  (),                        //               .bvalid
		.h2f_BREADY  (),                        //               .bready
		.h2f_ARID    (),                        //               .arid
		.h2f_ARADDR  (),                        //               .araddr
		.h2f_ARLEN   (),                        //               .arlen
		.h2f_ARSIZE  (),                        //               .arsize
		.h2f_ARBURST (),                        //               .arburst
		.h2f_ARLOCK  (),                        //               .arlock
		.h2f_ARCACHE (),                        //               .arcache
		.h2f_ARPROT  (),                        //               .arprot
		.h2f_ARVALID (),                        //               .arvalid
		.h2f_ARREADY (),                        //               .arready
		.h2f_RID     (),                        //               .rid
		.h2f_RDATA   (),                        //               .rdata
		.h2f_RRESP   (),                        //               .rresp
		.h2f_RLAST   (),                        //               .rlast
		.h2f_RVALID  (),                        //               .rvalid
		.h2f_RREADY  ()                         //               .rready
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (8),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (4),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (),                               //    s0.waitrequest
		.s0_readdata      (),                               //      .readdata
		.s0_readdatavalid (),                               //      .readdatavalid
		.s0_burstcount    (),                               //      .burstcount
		.s0_writedata     (),                               //      .writedata
		.s0_address       (),                               //      .address
		.s0_write         (),                               //      .write
		.s0_read          (),                               //      .read
		.s0_byteenable    (),                               //      .byteenable
		.s0_debugaccess   (),                               //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),         //      .address
		.m0_write         (mm_bridge_0_m0_write),           //      .write
		.m0_read          (mm_bridge_0_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),     //      .debugaccess
		.s0_response      (),                               // (terminated)
		.m0_response      (2'b00)                           // (terminated)
	);

	system_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pwm_input_0_export)                     // external_connection.export
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                               //                               clk_0_clk.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),        // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),            //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),             //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),             //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                   //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),               //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),          //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                  //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),              //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),            //                                        .debugaccess
		.pio_0_s1_address                              (mm_interconnect_0_pio_0_s1_address),    //                                pio_0_s1.address
		.pio_0_s1_write                                (mm_interconnect_0_pio_0_s1_write),      //                                        .write
		.pio_0_s1_readdata                             (mm_interconnect_0_pio_0_s1_readdata),   //                                        .readdata
		.pio_0_s1_writedata                            (mm_interconnect_0_pio_0_s1_writedata),  //                                        .writedata
		.pio_0_s1_chipselect                           (mm_interconnect_0_pio_0_s1_chipselect)  //                                        .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
